module gfg_verilog_Benchmark_testing100(I51,I59,I67,I75,I83,I91,I1403,I1417,I1445,I1470,I1526,I1540,I1565,I1621,I1635,I1660,I1702,I1716);
input I51,I59,I67,I75,I83,I91;
output I1403,I1417,I1445,I1470,I1526,I1540,I1565,I1621,I1635,I1660,I1702,I1716;
wire I51,I59,I67,I75,I83,I91,I99,I110,I124,I135,I146,I160,I174,I188,I202,I213,I224,I238,I249,I263,I277,I291,I305,I319,I333,I347,I361,I375,I389,I403,I414,I428,I442,I456,I470,I481,I495,I509,I520,I534,I548,I562,I576,I590,I604,I615,I629,I643,I657,I671,I685,I699,I713,I724,I738,I752,I766,I780,I794,I808,I819,I833,I847,I861,I875,I889,I903,I914,I928,I942,I956,I970,I984,I995,I1009,I1023,I1037,I1051,I1065,I1079,I1093,I1107,I1121,I1135,I1149,I1160,I1174,I1188,I1202,I1216,I1227,I1241,I1255,I1266,I1280,I1294,I1308,I1322,I1336,I1350,I1361,I1375,I1389,I1431,I1459,I1484,I1498,I1512,I1554,I1579,I1593,I1607,I1649,I1674,I1688;
buf I_6 (I99,I67);
nand I_7 (I110,I99,I51);
not I_8 (I124,I99);
buf I_9 (I135,I75);
nand I_10 (I146,I135,I124);
nand I_11 (I160,I146,I110);
nand I_12 (I174,I59,I83);
and I_13 (I188,I174,I51);
not I_14 (I202,I174);
not I_15 (I213,I91);
and I_16 (I224,I213,I202);
not I_17 (I238,I160);
nor I_18 (I249,I238,I99);
nor I_19 (I263,I124,I110);
nor I_20 (I277,I263,I160);
nor I_21 (I291,I277,I99);
nor I_22 (I305,I291,I124);
nor I_23 (I319,I238,I291);
nor I_24 (I333,I224,I188);
nor I_25 (I347,I333,I202);
nor I_26 (I361,I347,I213);
nor I_27 (I375,I333,I224);
nor I_28 (I389,I188,I202);
not I_29 (I403,I389);
nor I_30 (I414,I403,I361);
nor I_31 (I428,I389,I403);
nor I_32 (I442,I160,I135);
nor I_33 (I456,I442,I110);
not I_34 (I470,I160);
nor I_35 (I481,I470,I442);
nor I_36 (I495,I470,I135);
not I_37 (I509,I224);
nor I_38 (I520,I509,I188);
nor I_39 (I534,I202,I213);
nor I_40 (I548,I534,I224);
nor I_41 (I562,I548,I188);
nor I_42 (I576,I509,I562);
nor I_43 (I590,I534,I202);
not I_44 (I604,I319);
nor I_45 (I615,I305,I249);
nor I_46 (I629,I615,I277);
nor I_47 (I643,I629,I319);
nor I_48 (I657,I629,I643);
nor I_49 (I671,I604,I643);
nor I_50 (I685,I604,I305);
nor I_51 (I699,I685,I249);
not I_52 (I713,I428);
nor I_53 (I724,I713,I414);
nor I_54 (I738,I375,I333);
nor I_55 (I752,I738,I428);
nor I_56 (I766,I752,I414);
nor I_57 (I780,I766,I375);
nor I_58 (I794,I713,I766);
not I_59 (I808,I495);
nor I_60 (I819,I808,I481);
nor I_61 (I833,I456,I470);
nor I_62 (I847,I833,I495);
nor I_63 (I861,I847,I481);
nor I_64 (I875,I861,I456);
nor I_65 (I889,I808,I861);
not I_66 (I903,I590);
nor I_67 (I914,I903,I576);
and I_68 (I928,I520,I590);
nor I_69 (I942,I928,I576);
nor I_70 (I956,I942,I903);
nor I_71 (I970,I928,I942);
not I_72 (I984,I699);
nor I_73 (I995,I984,I671);
nor I_74 (I1009,I657,I629);
nor I_75 (I1023,I1009,I699);
nor I_76 (I1037,I1023,I671);
nor I_77 (I1051,I1037,I657);
nor I_78 (I1065,I984,I1037);
nor I_79 (I1079,I794,I780);
nor I_80 (I1093,I1079,I724);
nor I_81 (I1107,I1093,I738);
nor I_82 (I1121,I1079,I794);
nor I_83 (I1135,I780,I724);
not I_84 (I1149,I1135);
nor I_85 (I1160,I1149,I1107);
nor I_86 (I1174,I1135,I1149);
nor I_87 (I1188,I889,I875);
nor I_88 (I1202,I1188,I819);
not I_89 (I1216,I889);
nor I_90 (I1227,I1216,I1188);
nor I_91 (I1241,I1216,I875);
not I_92 (I1255,I970);
nor I_93 (I1266,I1255,I956);
nor I_94 (I1280,I914,I942);
nor I_95 (I1294,I1280,I970);
nor I_96 (I1308,I1294,I956);
nor I_97 (I1322,I1255,I1308);
nor I_98 (I1336,I1280,I914);
not I_99 (I1350,I1065);
nor I_100 (I1361,I1051,I995);
nor I_101 (I1375,I1361,I1023);
nor I_102 (I1389,I1375,I1065);
nor I_103 (I1403,I1375,I1389);
nor I_104 (I1417,I1350,I1389);
nor I_105 (I1431,I1350,I1051);
nor I_106 (I1445,I1431,I995);
not I_107 (I1459,I1174);
nor I_108 (I1470,I1459,I1160);
nor I_109 (I1484,I1121,I1079);
nor I_110 (I1498,I1484,I1174);
nor I_111 (I1512,I1498,I1160);
nor I_112 (I1526,I1512,I1121);
nor I_113 (I1540,I1459,I1512);
not I_114 (I1554,I1241);
nor I_115 (I1565,I1554,I1227);
nor I_116 (I1579,I1202,I1216);
nor I_117 (I1593,I1579,I1241);
nor I_118 (I1607,I1593,I1227);
nor I_119 (I1621,I1607,I1202);
nor I_120 (I1635,I1554,I1607);
not I_121 (I1649,I1336);
nor I_122 (I1660,I1649,I1322);
and I_123 (I1674,I1266,I1336);
nor I_124 (I1688,I1674,I1322);
nor I_125 (I1702,I1688,I1649);
nor I_126 (I1716,I1674,I1688);
endmodule


