module gfg_verilog_Benchmark_testing300(I51,I59,I67,I75,I83,I91,I3196,I3207,I3249,I3291,I3330,I3344,I3372,I3397,I3411,I3453,I3478,I3506,I3534,I3570,I3595,I3637,I3651,I3676,I3732,I3746,I3788,I3813,I3841,I3869,I3905,I3972,I3986,I3997,I4022,I4078,I4092);
input I51,I59,I67,I75,I83,I91;
output I3196,I3207,I3249,I3291,I3330,I3344,I3372,I3397,I3411,I3453,I3478,I3506,I3534,I3570,I3595,I3637,I3651,I3676,I3732,I3746,I3788,I3813,I3841,I3869,I3905,I3972,I3986,I3997,I4022,I4078,I4092;
wire I51,I59,I67,I75,I83,I91,I99,I110,I124,I135,I146,I160,I174,I188,I202,I213,I224,I238,I252,I266,I280,I294,I305,I319,I333,I344,I358,I372,I386,I400,I414,I428,I442,I453,I464,I478,I492,I506,I520,I531,I545,I559,I573,I587,I601,I615,I629,I643,I657,I668,I682,I696,I710,I724,I738,I749,I763,I774,I788,I802,I816,I830,I841,I855,I866,I880,I891,I905,I919,I933,I947,I961,I975,I989,I1003,I1017,I1031,I1042,I1056,I1067,I1081,I1092,I1106,I1120,I1134,I1148,I1162,I1176,I1187,I1201,I1212,I1223,I1237,I1251,I1262,I1273,I1287,I1301,I1315,I1329,I1343,I1357,I1371,I1385,I1396,I1410,I1424,I1438,I1452,I1463,I1477,I1491,I1505,I1519,I1533,I1544,I1558,I1572,I1586,I1600,I1614,I1625,I1636,I1650,I1661,I1675,I1689,I1703,I1717,I1731,I1742,I1756,I1770,I1784,I1798,I1812,I1826,I1840,I1854,I1868,I1879,I1893,I1907,I1921,I1935,I1949,I1960,I1971,I1985,I1999,I2013,I2027,I2038,I2052,I2063,I2077,I2088,I2102,I2116,I2130,I2144,I2158,I2172,I2186,I2200,I2214,I2228,I2239,I2253,I2267,I2278,I2292,I2306,I2320,I2334,I2348,I2362,I2376,I2387,I2398,I2412,I2426,I2440,I2454,I2465,I2479,I2493,I2507,I2521,I2535,I2549,I2563,I2577,I2591,I2602,I2616,I2630,I2644,I2658,I2672,I2683,I2697,I2708,I2722,I2736,I2750,I2764,I2775,I2789,I2800,I2814,I2825,I2839,I2853,I2867,I2881,I2895,I2909,I2923,I2937,I2951,I2965,I2976,I2990,I3001,I3015,I3026,I3040,I3054,I3068,I3082,I3096,I3110,I3121,I3135,I3146,I3157,I3171,I3185,I3221,I3235,I3263,I3277,I3305,I3319,I3358,I3386,I3425,I3439,I3467,I3492,I3520,I3548,I3559,I3584,I3609,I3623,I3665,I3690,I3704,I3718,I3760,I3774,I3802,I3827,I3855,I3883,I3894,I3919,I3933,I3947,I3961,I4011,I4036,I4050,I4064;
buf I_6 (I99,I67);
nand I_7 (I110,I99,I83);
not I_8 (I124,I99);
buf I_9 (I135,I59);
nand I_10 (I146,I135,I124);
nand I_11 (I160,I146,I110);
nand I_12 (I174,I51,I91);
and I_13 (I188,I174,I75);
not I_14 (I202,I174);
not I_15 (I213,I67);
and I_16 (I224,I213,I202);
and I_17 (I238,I160,I135);
nor I_18 (I252,I238,I146);
nor I_19 (I266,I238,I252);
and I_20 (I280,I160,I135);
not I_21 (I294,I280);
nor I_22 (I305,I294,I252);
nor I_23 (I319,I280,I294);
not I_24 (I333,I224);
nor I_25 (I344,I188,I213);
nor I_26 (I358,I344,I202);
nor I_27 (I372,I358,I224);
nor I_28 (I386,I358,I372);
nor I_29 (I400,I333,I372);
nor I_30 (I414,I333,I188);
nor I_31 (I428,I414,I213);
not I_32 (I442,I160);
not I_33 (I453,I442);
nor I_34 (I464,I442,I135);
and I_35 (I478,I124,I160);
nor I_36 (I492,I478,I135);
nor I_37 (I506,I492,I442);
not I_38 (I520,I160);
nor I_39 (I531,I520,I146);
and I_40 (I545,I110,I160);
nor I_41 (I559,I545,I146);
nor I_42 (I573,I559,I520);
nor I_43 (I587,I545,I559);
and I_44 (I601,I224,I188);
nor I_45 (I615,I601,I213);
nor I_46 (I629,I601,I615);
and I_47 (I643,I224,I188);
not I_48 (I657,I643);
nor I_49 (I668,I657,I615);
nor I_50 (I682,I643,I657);
and I_51 (I696,I160,I135);
nor I_52 (I710,I696,I99);
and I_53 (I724,I160,I135);
not I_54 (I738,I724);
nor I_55 (I749,I738,I710);
not I_56 (I763,I738);
nor I_57 (I774,I724,I738);
and I_58 (I788,I160,I135);
nor I_59 (I802,I788,I99);
and I_60 (I816,I160,I135);
not I_61 (I830,I816);
nor I_62 (I841,I830,I802);
not I_63 (I855,I830);
nor I_64 (I866,I816,I830);
not I_65 (I880,I160);
nor I_66 (I891,I124,I110);
nor I_67 (I905,I891,I99);
nor I_68 (I919,I905,I160);
nor I_69 (I933,I905,I919);
nor I_70 (I947,I880,I919);
nor I_71 (I961,I880,I124);
nor I_72 (I975,I961,I110);
nor I_73 (I989,I160,I99);
nor I_74 (I1003,I989,I124);
nor I_75 (I1017,I160,I99);
not I_76 (I1031,I1017);
nor I_77 (I1042,I1031,I1003);
not I_78 (I1056,I1031);
nor I_79 (I1067,I1017,I1031);
not I_80 (I1081,I224);
nor I_81 (I1092,I1081,I188);
nor I_82 (I1106,I202,I174);
nor I_83 (I1120,I1106,I224);
nor I_84 (I1134,I1120,I188);
nor I_85 (I1148,I1134,I202);
nor I_86 (I1162,I1081,I1134);
buf I_87 (I1176,I224);
nand I_88 (I1187,I1176,I188);
not I_89 (I1201,I1176);
buf I_90 (I1212,I224);
nand I_91 (I1223,I1212,I1201);
nand I_92 (I1237,I1223,I1187);
not I_93 (I1251,I319);
not I_94 (I1262,I1251);
nor I_95 (I1273,I1251,I305);
and I_96 (I1287,I266,I319);
nor I_97 (I1301,I1287,I305);
nor I_98 (I1315,I1301,I1251);
and I_99 (I1329,I975,I947);
nor I_100 (I1343,I1329,I933);
nor I_101 (I1357,I1329,I1343);
and I_102 (I1371,I975,I947);
not I_103 (I1385,I1371);
nor I_104 (I1396,I1385,I1343);
nor I_105 (I1410,I1371,I1385);
nor I_106 (I1424,I506,I464);
nor I_107 (I1438,I1424,I453);
not I_108 (I1452,I506);
nor I_109 (I1463,I1452,I1424);
nor I_110 (I1477,I1452,I464);
nor I_111 (I1491,I587,I573);
nor I_112 (I1505,I1491,I531);
nor I_113 (I1519,I1505,I545);
not I_114 (I1533,I587);
nor I_115 (I1544,I1533,I1505);
nor I_116 (I1558,I1533,I573);
nor I_117 (I1572,I1558,I531);
nand I_118 (I1586,I682,I668);
and I_119 (I1600,I1586,I629);
not I_120 (I1614,I1586);
not I_121 (I1625,I682);
and I_122 (I1636,I1625,I1614);
not I_123 (I1650,I866);
nor I_124 (I1661,I1650,I855);
and I_125 (I1675,I841,I866);
nor I_126 (I1689,I1675,I855);
nor I_127 (I1703,I1689,I1650);
nor I_128 (I1717,I1675,I1689);
not I_129 (I1731,I774);
nor I_130 (I1742,I1731,I763);
nor I_131 (I1756,I749,I710);
nor I_132 (I1770,I1756,I774);
nor I_133 (I1784,I1770,I763);
nor I_134 (I1798,I1784,I749);
nor I_135 (I1812,I1731,I1784);
nor I_136 (I1826,I428,I400);
nor I_137 (I1840,I1826,I386);
nor I_138 (I1854,I1840,I372);
not I_139 (I1868,I428);
nor I_140 (I1879,I1868,I1840);
nor I_141 (I1893,I1868,I400);
nor I_142 (I1907,I1893,I386);
nand I_143 (I1921,I1067,I1056);
and I_144 (I1935,I1921,I1042);
not I_145 (I1949,I1921);
not I_146 (I1960,I1067);
and I_147 (I1971,I1960,I1949);
nor I_148 (I1985,I1162,I1148);
nor I_149 (I1999,I1985,I1092);
nor I_150 (I2013,I1162,I1148);
not I_151 (I2027,I2013);
nor I_152 (I2038,I2027,I1999);
not I_153 (I2052,I2027);
nor I_154 (I2063,I2013,I2027);
not I_155 (I2077,I1237);
nor I_156 (I2088,I2077,I1187);
nor I_157 (I2102,I1176,I1212);
nor I_158 (I2116,I2102,I1237);
nor I_159 (I2130,I2116,I1187);
nor I_160 (I2144,I2077,I2130);
nor I_161 (I2158,I2102,I1176);
and I_162 (I2172,I1315,I1273);
nor I_163 (I2186,I2172,I1262);
nor I_164 (I2200,I2172,I2186);
and I_165 (I2214,I1315,I1273);
not I_166 (I2228,I2214);
nor I_167 (I2239,I2228,I2186);
nor I_168 (I2253,I2214,I2228);
not I_169 (I2267,I1410);
nor I_170 (I2278,I1396,I1357);
nor I_171 (I2292,I2278,I1343);
nor I_172 (I2306,I2292,I1410);
nor I_173 (I2320,I2292,I2306);
nor I_174 (I2334,I2267,I2306);
nor I_175 (I2348,I2267,I1396);
nor I_176 (I2362,I2348,I1357);
not I_177 (I2376,I1477);
not I_178 (I2387,I2376);
nor I_179 (I2398,I2376,I1463);
and I_180 (I2412,I1438,I1477);
nor I_181 (I2426,I2412,I1463);
nor I_182 (I2440,I2426,I2376);
not I_183 (I2454,I1572);
nor I_184 (I2465,I2454,I1544);
and I_185 (I2479,I1519,I1572);
nor I_186 (I2493,I2479,I1544);
nor I_187 (I2507,I2493,I2454);
nor I_188 (I2521,I2479,I2493);
and I_189 (I2535,I1636,I1600);
nor I_190 (I2549,I2535,I1625);
nor I_191 (I2563,I2535,I2549);
and I_192 (I2577,I1636,I1600);
not I_193 (I2591,I2577);
nor I_194 (I2602,I2591,I2549);
nor I_195 (I2616,I2577,I2591);
and I_196 (I2630,I1717,I1703);
nor I_197 (I2644,I2630,I1661);
and I_198 (I2658,I1717,I1703);
not I_199 (I2672,I2658);
nor I_200 (I2683,I2672,I2644);
not I_201 (I2697,I2672);
nor I_202 (I2708,I2658,I2672);
and I_203 (I2722,I1812,I1798);
nor I_204 (I2736,I2722,I1742);
and I_205 (I2750,I1812,I1798);
not I_206 (I2764,I2750);
nor I_207 (I2775,I2764,I2736);
not I_208 (I2789,I2764);
nor I_209 (I2800,I2750,I2764);
not I_210 (I2814,I1907);
nor I_211 (I2825,I1879,I1854);
nor I_212 (I2839,I2825,I1893);
nor I_213 (I2853,I2839,I1907);
nor I_214 (I2867,I2839,I2853);
nor I_215 (I2881,I2814,I2853);
nor I_216 (I2895,I2814,I1879);
nor I_217 (I2909,I2895,I1854);
nor I_218 (I2923,I1971,I1935);
nor I_219 (I2937,I2923,I1921);
nor I_220 (I2951,I1971,I1935);
not I_221 (I2965,I2951);
nor I_222 (I2976,I2965,I2937);
not I_223 (I2990,I2965);
nor I_224 (I3001,I2951,I2965);
not I_225 (I3015,I2063);
nor I_226 (I3026,I3015,I2052);
nor I_227 (I3040,I2038,I1999);
nor I_228 (I3054,I3040,I2063);
nor I_229 (I3068,I3054,I2052);
nor I_230 (I3082,I3068,I2038);
nor I_231 (I3096,I3015,I3068);
buf I_232 (I3110,I2158);
nand I_233 (I3121,I3110,I2144);
not I_234 (I3135,I3110);
buf I_235 (I3146,I2088);
nand I_236 (I3157,I3146,I3135);
nand I_237 (I3171,I3157,I3121);
not I_238 (I3185,I2616);
not I_239 (I3196,I3185);
nor I_240 (I3207,I3185,I2602);
and I_241 (I3221,I2563,I2616);
nor I_242 (I3235,I3221,I2602);
nor I_243 (I3249,I3235,I3185);
and I_244 (I3263,I2362,I2334);
nor I_245 (I3277,I3263,I2320);
nor I_246 (I3291,I3263,I3277);
and I_247 (I3305,I2362,I2334);
not I_248 (I3319,I3305);
nor I_249 (I3330,I3319,I3277);
nor I_250 (I3344,I3305,I3319);
nor I_251 (I3358,I2440,I2398);
nor I_252 (I3372,I3358,I2387);
not I_253 (I3386,I2440);
nor I_254 (I3397,I3386,I3358);
nor I_255 (I3411,I3386,I2398);
nor I_256 (I3425,I2521,I2507);
nor I_257 (I3439,I3425,I2465);
nor I_258 (I3453,I3439,I2479);
not I_259 (I3467,I2521);
nor I_260 (I3478,I3467,I3439);
nor I_261 (I3492,I3467,I2507);
nor I_262 (I3506,I3492,I2465);
nand I_263 (I3520,I2253,I2239);
and I_264 (I3534,I3520,I2200);
not I_265 (I3548,I3520);
not I_266 (I3559,I2253);
and I_267 (I3570,I3559,I3548);
not I_268 (I3584,I2708);
nor I_269 (I3595,I3584,I2697);
and I_270 (I3609,I2683,I2708);
nor I_271 (I3623,I3609,I2697);
nor I_272 (I3637,I3623,I3584);
nor I_273 (I3651,I3609,I3623);
not I_274 (I3665,I2800);
nor I_275 (I3676,I3665,I2789);
nor I_276 (I3690,I2775,I2736);
nor I_277 (I3704,I3690,I2800);
nor I_278 (I3718,I3704,I2789);
nor I_279 (I3732,I3718,I2775);
nor I_280 (I3746,I3665,I3718);
nor I_281 (I3760,I2909,I2881);
nor I_282 (I3774,I3760,I2867);
nor I_283 (I3788,I3774,I2853);
not I_284 (I3802,I2909);
nor I_285 (I3813,I3802,I3774);
nor I_286 (I3827,I3802,I2881);
nor I_287 (I3841,I3827,I2867);
nand I_288 (I3855,I3001,I2990);
and I_289 (I3869,I3855,I2976);
not I_290 (I3883,I3855);
not I_291 (I3894,I3001);
and I_292 (I3905,I3894,I3883);
nor I_293 (I3919,I3096,I3082);
nor I_294 (I3933,I3919,I3026);
nor I_295 (I3947,I3096,I3082);
not I_296 (I3961,I3947);
nor I_297 (I3972,I3961,I3933);
not I_298 (I3986,I3961);
nor I_299 (I3997,I3947,I3961);
not I_300 (I4011,I3171);
nor I_301 (I4022,I4011,I3121);
nor I_302 (I4036,I3110,I3146);
nor I_303 (I4050,I4036,I3171);
nor I_304 (I4064,I4050,I3121);
nor I_305 (I4078,I4011,I4064);
nor I_306 (I4092,I4036,I3110);
endmodule


